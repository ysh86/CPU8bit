module SW (
  input  logic nIN,
  output logic nOUT
);

  assign nOUT = nIN;

endmodule
